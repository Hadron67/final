module TLB #(
    parameter ENTRY_ADDR_WIDTH = 3;
) (
    
);

endmodule // TLB