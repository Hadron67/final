module spi_tb();
    
    SPIMaster spi();
endmodule