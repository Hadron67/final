interface CPUControl;
    wire aluSrcA;
    wire aluSrcB;
    wire aluOptr;
    wire aluOverflow;
    wire regDest;
    wire extOp;
    wire writeReg;
    wire writeRegSrc;
    wire writeMem;
    wire readMem;
    wire jmp;
    wire branch;
    wire branchCond;
endinterface