`include "DataBus.vh"

module CachTop(
        
);

endmodule // CachTop