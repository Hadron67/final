module mmu_tb();
    MMU uut ();
endmodule // mmu_tb